module conspiracion;
endmodule
