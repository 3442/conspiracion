`ifndef CORE_PSR_SV
`define CORE_PSR_SV

typedef struct packed
{
	logic n, z, c, v;
} psr_flags;

`endif
