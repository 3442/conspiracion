`ifndef CORE_CP15_MAP_SV
`define CORE_CP15_MAP_SV

`define CP15_CRN_CPUID     4'd0
`define CP15_CRN_SYSCFG    4'd1
`define CP15_CRN_TTBR      4'd2
`define CP15_CRN_DOMAIN    4'd3
`define CP15_CRN_FSR       4'd5
`define CP15_CRN_FAR       4'd6
`define CP15_CRN_CACHE     4'd7
`define CP15_CRN_TLB       4'd8
`define CP15_CRN_CACHE_LCK 4'd9
`define CP15_CRN_TLB_LCK   4'd10
`define CP15_CRN_DMA       4'd11
`define CP15_CRN_PID       4'd13

`endif
