`ifndef CONFIG_SV
`define CONFIG_SV

`define CONFIG_CPUS  1
`define CONFIG_CACHE 1

`endif
