`include "core/uarch.sv"

module core_cp15_tlb
(
	input  logic     clk,
	                 rst_n,

	input  logic     load,
	                 transfer,
	input  word      write
);

	//TODO

endmodule
