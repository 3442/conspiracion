`include "core/mmu/format.sv"
`include "core/uarch.sv"

module core_mmu
(
	input  logic      clk,
	                  rst_n,

	input  logic      mmu_enable /*verilator public*/,
	input  mmu_base   mmu_ttbr /*verilator public*/,

	input  logic      bus_ready,
	input  word       bus_data_rd,
	                  data_data_wr,
	input  ptr        insn_addr,
	                  data_addr,
	input  logic      insn_start,
	                  data_start,
	                  data_write,
	input  logic[3:0] data_data_be,

	output word       bus_data_wr,
	output logic[3:0] bus_data_be,
	output ptr        bus_addr,
	output logic      bus_start,
	                  bus_write,
	                  insn_ready,
	                  data_ready,
	                  data_fault,
	output word       insn_data_rd,
	                  data_data_rd,

	output logic      fault_register,
	output ptr        fault_addr
);

	ptr iphys_addr, dphys_addr;
	word iphys_data_rd, dphys_data_rd, dphys_data_wr;
	logic iphys_start, dphys_start, iphys_ready, dphys_ready, dphys_write;
	logic[3:0] dphys_data_be;

	assign fault_register = data_fault;

	core_mmu_pagewalk iwalk
	(
		.core_addr(insn_addr),
		.core_start(insn_start),
		.core_write(0),
		.core_ready(insn_ready),
		.core_fault(),
		.core_data_wr(0),
		.core_data_be(0),
		.core_data_rd(insn_data_rd),
		.core_fault_addr(),

		.bus_addr(iphys_addr),
		.bus_start(iphys_start),
		.bus_write(),
		.bus_ready(iphys_ready),
		.bus_data_wr(),
		.bus_data_be(),
		.bus_data_rd(iphys_data_rd),

		.*
	);

	core_mmu_pagewalk dwalk
	(
		.core_addr(data_addr),
		.core_start(data_start),
		.core_write(data_write),
		.core_ready(data_ready),
		.core_fault(data_fault),
		.core_data_wr(data_data_wr),
		.core_data_be(data_data_be),
		.core_data_rd(data_data_rd),
		.core_fault_addr(fault_addr),

		.bus_addr(dphys_addr),
		.bus_start(dphys_start),
		.bus_write(dphys_write),
		.bus_ready(dphys_ready),
		.bus_data_wr(dphys_data_wr),
		.bus_data_be(dphys_data_be),
		.bus_data_rd(dphys_data_rd),

		.*
	);

	core_mmu_arbiter arbiter
	(
		.insn_addr(iphys_addr),
		.insn_start(iphys_start),
		.insn_ready(iphys_ready),
		.insn_data_rd(iphys_data_rd),

		.data_addr(dphys_addr),
		.data_start(dphys_start),
		.data_write(dphys_write),
		.data_ready(dphys_ready),
		.data_data_wr(dphys_data_wr),
		.data_data_be(dphys_data_be),
		.data_data_rd(dphys_data_rd),

		.*
	);

endmodule
