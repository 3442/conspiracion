`include "core/uarch.sv"

module core_cp15_cache
(
	input  logic     clk,
	                 rst_n,

	input  logic     load,
	                 transfer,
	input  word      write
);

	//TODO

endmodule
