`ifndef CONFIG_SV
`define CONFIG_SV

`define CONFIG_CPUS         4
`define CONFIG_CACHE        1
`define CONFIG_PERF_MONITOR 1

`endif
